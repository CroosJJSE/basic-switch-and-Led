`timescale 1ns / 1ps

module top(
    input switch,
    output led
    );
    assign led = switch ;
endmodule
